`include "Arabi.Sina.400243058.Problem1.v"

module Q1_tb();
    reg A, B, C, D;
    wire out;
    f f(out, A, B, C, D);

initial begin
    A = 0;
    B = 0;
    C = 0;
    D = 0;
#20;
    A = 0;
    B = 0;
    C = 0;
    D = 1;
#20;
    A = 0;
    B = 0;
    C = 1;
    D = 0;
#20;
    A = 0;
    B = 0;
    C = 1;
    D = 1;
#20;
    A = 0;
    B = 1;
    C = 0;
    D = 0;
#20;
    A = 0;
    B = 1;
    C = 0;
    D = 1;
#20;
    A = 0;
    B = 1;
    C = 1;
    D = 0;
#20;
    A = 0;
    B = 1;
    C = 1;
    D = 1;
#20;
    A = 1;
    B = 0;
    C = 0;
    D = 0;
#20;
    A = 1;
    B = 0;
    C = 0;
    D = 1;
#20;
    A = 1;
    B = 0;
    C = 1;
    D = 0;
#20;
    A = 1;
    B = 0;
    C = 1;
    D = 1;
#20;
    A = 1;
    B = 1;
    C = 0;
    D = 0;
#20;
    A = 1;
    B = 1;
    C = 0;
    D = 1;
#20;
    A = 1;
    B = 1;
    C = 1;
    D = 0;
#20;
    A = 1;
    B = 1;
    C = 1;
    D = 1;
#20;
end

endmodule
